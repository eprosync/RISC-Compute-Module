// FPU - Floating Point Unit
// This is a LOT more complicated than an ALU
// Since now we have to deal with IEEE 754
// 32 - 1 bit (sign) | 8 bits (exponent) | 23 bits (mantissa)
// 64 - 1 bit (sign) | 11 bits (exponent) | 52 bits (mantissa)

module FPU ()

endmodule